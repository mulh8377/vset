module main
fn main () {}
